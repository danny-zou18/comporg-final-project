module arch;

    // Define signals for testbench inputs and outputs
    reg clk;
    reg reset;
    // Define other necessary testbench signals
    
    // Instantiate the CPU module
    CPU dut (
        .clk(clk),
        .reset(reset),
        // Connect other inputs and outputs
        // Example:
        .address_bus(...), // Connect appropriate signals from testbench
        .data_bus_in(...), // Connect appropriate signals from testbench
        .data_bus_out(...) // Connect appropriate signals from testbench
    );

    // Clock generation
    always #5 clk = ~clk;  // Example: Generate a clock signal

    // Initial stimulus
    initial begin
        clk = 0;
        reset = 1;  // Apply reset initially
        // Apply other initial stimuli
        
        #50 reset = 0;  // Deassert reset after some time
        
        // Add more testbench stimulus and checks here
        // For example: apply inputs and monitor outputs
        
        #1000 $finish;  // End simulation after certain time
    end

endmodule
